// Greg Stitt
// Wes Piard
// University of Florida

`ifndef _AXI4_STREAM_IF_
`define _AXI4_STREAM_IF_

interface axi4_stream_if #(
    parameter int DATA_WIDTH = 64,
    parameter int ID_WIDTH   = 0,
    parameter int DEST_WIDTH = 0,
    parameter int USER_WIDTH = 0
) (
    input logic aclk,
    input logic aresetn
);
    logic tvalid;
    logic tready;
    logic [DATA_WIDTH-1:0] tdata;
    logic [DATA_WIDTH/8-1:0] tstrb;
    logic [DATA_WIDTH/8-1:0] tkeep;
    logic tlast;
    logic [ID_WIDTH-1:0] tid;
    logic [DEST_WIDTH-1:0] tdest;
    logic [USER_WIDTH-1:0] tuser;

    // ===================================
    // MODPORTS
    // ===================================

    modport Source(input aclk, aresetn, input tready, output tvalid, tdata, tstrb, tkeep, tlast, tuser, tid, tdest, import clear_source_outputs);

    modport Sink(input aclk, aresetn, input tvalid, tdata, tstrb, tkeep, tlast, tuser, tid, tdest, output tready, import clear_sink_outputs);

    // AXI requires byte-aligned data widths, so confirm compliance here.
    initial begin
        if (DATA_WIDTH % 8 != 0) $fatal(1, $sformatf("AXI DATA_WIDTH=%0d is not byte aligned", DATA_WIDTH));
    end

    // Validate required properties of AXI: once tvalid is asserted, it must remain asserted until
    // tready is asserted.
    assert property (@(posedge aclk) disable iff (!aresetn) $fell(tvalid) |-> $past(tready, 1))
    else $error("tvalid must be asserted continuously until tready is asserted.");

endinterface

`endif
